module m21_32_bit(Y, D0, D1, S);
input S;
input [31:0]D0,D1;
output [31:0]Y;

m21 q0(Y[0], D0[0], D1[0],S);
m21 q1(Y[1], D0[1], D1[1],S);
m21 q2(Y[2], D0[2], D1[2],S);
m21 q3(Y[3], D0[3], D1[3],S);
m21 q4(Y[4], D0[4], D1[4],S);
m21 q5(Y[5], D0[5], D1[5],S);
m21 q6(Y[6], D0[6], D1[6],S);
m21 q7(Y[7], D0[7], D1[7],S);
m21 q8(Y[8], D0[8], D1[8],S);
m21 q9(Y[9], D0[9], D1[9],S);
m21 q10(Y[10], D0[10], D1[10],S);
m21 q11(Y[11], D0[11], D1[11],S);
m21 q12(Y[12], D0[12], D1[12], S);
m21 q13(Y[13], D0[13], D1[13], S);
m21 q14(Y[14], D0[14], D1[14], S);
m21 q15(Y[15], D0[15], D1[15], S);
m21 q16(Y[16], D0[16], D1[16], S);
m21 q17(Y[17], D0[17], D1[17], S);
m21 q18(Y[18], D0[18], D1[18], S);
m21 q19(Y[19], D0[19], D1[19], S);
m21 q20(Y[20], D0[20], D1[20], S);
m21 q21(Y[21], D0[21], D1[21], S);
m21 q22(Y[22], D0[22], D1[22], S);
m21 q23(Y[23], D0[23], D1[23], S);
m21 q24(Y[24], D0[24], D1[24], S);
m21 q25(Y[25], D0[25], D1[25], S);
m21 q26(Y[26], D0[26], D1[26], S);
m21 q27(Y[27], D0[27], D1[27], S);
m21 q28(Y[28], D0[28], D1[28], S);
m21 q29(Y[29], D0[29], D1[29], S);
m21 q30(Y[30], D0[30], D1[30], S);
m21 q31(Y[31], D0[31], D1[31], S);
endmodule