module Myps();
Instruction_Memory(pc,instructionn);

endmodule